`default_nettype wire



















